library verilog;
use verilog.vl_types.all;
entity Ula_1bit_vlg_vec_tst is
end Ula_1bit_vlg_vec_tst;
