library verilog;
use verilog.vl_types.all;
entity Full_Adder_1_bit_vlg_vec_tst is
end Full_Adder_1_bit_vlg_vec_tst;
